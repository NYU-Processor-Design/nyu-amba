/**
  @brief APB Bridge implementation

  @note See https://developer.arm.com/documentation/ihi0011/a/AMBA-APB/APB-bridge/Interface-diagram
*/
module Bridge (
  AHBCommon_if.subordinate sub,
  APBCommon_if.bridge bridge
);
  // Interface the two modports here

endmodule
