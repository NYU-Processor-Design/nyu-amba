/**
  @brief Subordinate to interface witht he memory controller

  @note See https://github.com/NYU-Processor-Design/nyu-mem
*/

module SubMemCtrl(
  AHBCommon_if.subordinate sub,
  MemCommon_if.memCtrl mem
);
  // General subordinate logic follows

endmodule
